module hcms_serial (
    input CLK_i
);
    


endmodule