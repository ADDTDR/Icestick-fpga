module top (
    input PMOD_4,
    input PMOD_3,
    output D1,
    output D2
);
    assign D1 = PMOD_4;
    assign D2 = PMOD_3;

endmodule